CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 40 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 6 110 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100626 0
0
6 Title:
5 Name:
0
0
0
10
6 74LS48
188 819 443 0 14 29
0 11 12 14 13 26 27 5 6 7
2 8 9 10 28
0
0 0 4832 0
6 74LS48
-20 59 22 67
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5130 0 0
2
43530.5 9
0
6 74112~
219 325 370 0 7 32
0 4 4 3 4 4 25 13
0
0 0 4704 0
5 74112
-72 -24 -37 -16
3 FFA
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
391 0 0
2
43530.5 8
0
6 74112~
219 451 370 0 7 32
0 4 13 3 13 4 24 14
0
0 0 4704 0
5 74112
-71 -23 -36 -15
3 FFB
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3124 0 0
2
43530.5 7
0
6 74112~
219 577 370 0 7 32
0 4 16 3 16 4 23 12
0
0 0 4704 0
5 74112
-72 -23 -37 -15
3 FFC
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3421 0 0
2
43530.5 6
0
6 74112~
219 703 370 0 7 32
0 4 15 3 15 4 22 11
0
0 0 4704 0
5 74112
-72 -22 -37 -14
3 FFD
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8157 0 0
2
43530.5 5
0
9 2-In AND~
219 522 254 0 3 22
0 13 14 16
0
0 0 608 0
6 74LS08
-24 21 18 29
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43530.5 4
0
9 2-In AND~
219 649 253 0 3 22
0 16 12 15
0
0 0 608 0
6 74LS08
-25 22 17 30
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
43530.5 3
0
9 CC 7-Seg~
183 918 332 0 18 19
10 10 9 8 2 7 6 5 20 21
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
6 BLUECC
-76 -3 -34 5
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7361 0 0
2
43530.5 2
0
7 Pulser~
4 138 346 0 10 12
0 17 18 3 19 0 0 5 5 6
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4747 0 0
2
43530.5 1
0
2 +V
167 325 264 0 1 3
0 4
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
43530.5 0
0
35
10 4 2 0 0 16 0 1 8 0 0 3
851 434
915 434
915 368
3 0 3 0 0 16 0 2 0 0 10 2
295 343
295 399
2 1 4 0 0 16 0 2 10 0 0 3
301 334
301 273
325 273
4 2 4 0 0 16 0 2 2 0 0 2
301 352
301 334
0 0 4 0 0 16 0 0 0 6 13 2
371 307
371 382
1 1 4 0 0 16 0 2 3 0 0 2
325 307
451 307
1 1 4 0 0 16 0 10 2 0 0 2
325 273
325 307
3 0 3 0 0 16 0 3 0 0 10 2
421 343
421 399
3 0 3 0 0 16 0 4 0 0 10 2
547 343
547 399
3 3 3 0 0 16 0 9 5 0 0 5
162 337
214 337
214 399
673 399
673 343
5 5 4 0 0 16 0 4 5 0 0 2
577 382
703 382
5 5 4 0 0 16 0 3 4 0 0 2
451 382
577 382
5 5 4 0 0 16 0 2 3 0 0 2
325 382
451 382
7 7 5 0 0 16 0 1 8 0 0 3
851 407
933 407
933 368
8 6 6 0 0 16 0 1 8 0 0 3
851 416
927 416
927 368
9 5 7 0 0 16 0 1 8 0 0 3
851 425
921 425
921 368
11 3 8 0 0 16 0 1 8 0 0 3
851 443
909 443
909 368
12 2 9 0 0 16 0 1 8 0 0 3
851 452
903 452
903 368
13 1 10 0 0 16 0 1 8 0 0 3
851 461
897 461
897 368
1 7 11 0 0 16 0 1 5 0 0 3
787 407
727 407
727 334
7 2 12 0 0 16 0 4 1 0 0 3
601 334
601 416
787 416
7 4 13 0 0 16 0 2 1 0 0 3
349 334
349 434
787 434
3 7 14 0 0 16 0 1 3 0 0 3
787 425
475 425
475 334
2 3 15 0 0 16 0 5 7 0 0 3
679 334
679 253
670 253
2 7 12 0 0 16 0 7 4 0 0 3
625 262
625 334
601 334
3 1 16 0 0 16 0 6 7 0 0 4
543 254
612 254
612 244
625 244
2 3 16 0 0 16 0 4 6 0 0 3
553 334
553 254
543 254
2 1 13 0 0 16 0 3 6 0 0 3
427 334
427 245
498 245
7 2 14 0 0 16 0 3 6 0 0 3
475 334
475 263
498 263
7 2 13 0 0 16 0 2 3 0 0 2
349 334
427 334
2 4 15 0 0 16 0 5 5 0 0 2
679 334
679 352
2 4 16 0 0 16 0 4 4 0 0 2
553 334
553 352
2 4 13 0 0 16 0 3 3 0 0 2
427 334
427 352
1 1 4 0 0 16 0 4 5 0 0 2
577 307
703 307
1 1 4 0 0 16 0 3 4 0 0 2
451 307
577 307
2
-27 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 24
16 60 412 113
25 67 402 102
24 Derek G. Apit BSCpE - 1B
-32 0 0 0 700 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 35
151 137 1043 199
164 145 1029 187
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
